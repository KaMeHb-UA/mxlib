module mxlib

fn test_init() ? {
	init('https', 'matrix.org', 443)?
}
